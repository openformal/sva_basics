/*md
# Description
This testbench explains concurrancy in concurrent sequences.

# DUT
This testbench uses a round robin arbiter as a context for introducing the
concepts. The dut design file is -
[sva_basics/design/src/rr_arbiter.sv](https://github.com/openformal/sva_basics/blob/master/design/docs/rr_arbiter.md)

*/

//sv+
module concurrency_tb();

  logic clock;
  logic reset;

  parameter CLIENTS = 32;

  logic [CLIENTS-1:0] request;
  logic [CLIENTS-1:0] grant;

//md In this testbench stall is disabled
  wire stall = 1'b0;

  rr_arbiter #(.CLIENTS(32)) dut (
                  .request (request),
                  .grant   (grant),
                  .stall   (stall),
                  .clock   (clock),
                  .reset   (reset));

/*md
# Overview
Concurrent SVAs are evaluated every clock cycle. Each one is a separate thread
that spans one or multiple clock cycles.

Consider the cover property below.
*/
  sequence gnt4_in_31_cycles_S;
    request[4] ##[0:31] grant[4];
  endsequence;

  gnt4_in_31_cycles_C: cover property (
    @(posedge clock) (gnt4_in_31_cycles_S)
  );

/*md
Now consider a scenario where request[4] is asserted at cycle *n*
and grant arrives at cycle *n+10*.
Between the cycle *n* to *n+10* the cover will start a new thread 11 times,
because concurrent assetions start a thread every cycle.
On cycle *n+10* 11 covers will finish, ranging from 0-10 cycles long.
/*md

# Concurrency wrt formal verification

The above example is more simulation centric as the scenario is preknown.
In formal verification the scenarios are generated by the tool. It is still
important to pay attention to concurrency.

Consider a verion of an arbiter that has requests and grants as single cycle
pulses. This arbiter allows upto 4 outstanding requests per requestor. If not
carefully code a single grant will satisfy multiple requests in the
testbench.
*/
/*md
# Avoiding muliple concurrent multicycle threads
In the dut above, the arbiter requires the request to be held high till
grant is received. Below is another way of writing the cover property above.
*$rose* for a bit is true at when it goes it is sampled 0 the previous cycle
and 1 in the current cycle.
This cover will also start 11 instances. But 10 of those 11 instances will
finish the cycle they start because of the use of *$rose*. At the *n+11* cycle
there will be only one match, and it will be for the cover that started at
cycle *n*
*/

  gnt4_in_31_cycles_C1: cover property (
    @(posedge clock) $rose(request[4]) ##[0:31] grant[4]
  );

endmodule
//sv-
